/*
设计一个能够有多种工作模式控制的8个灯亮灭的电路。
工作模式1：按照从左到右的方向，依次点亮每一盏灯，然后依次熄灭每一盏灯；
工作模式2：分成两组灯，前四个灯为1组，后四个为2组，1组灯按从左到右依次点亮，同时2组灯按从右到左依次点亮，然后两组灯按各自点亮的顺序依次熄灭；
工作模式3：用11110000作为一组灯的序列，按照该顺序完成8盏灯亮灭：即首先灯1亮，然后灯2亮，然后灯3亮，然后灯4亮，然后灯5不亮，然后灯6不亮，然后灯7不亮，然后灯8不亮，然后八个灯同时变成亮，亮，亮，亮，不亮，不亮，不亮，不亮，并保持下去。
工作模式4：自行设计一个模式控制8个灯亮灭。要求和前三个工作模式不同。

要求每种工作模式重复两次，并在2分钟内完成所有工作模式。
输入信号： 选择信号[1:0]S, 时钟信号clk, 复位信号reset
输出信号： 跑马灯亮灭信号[7:0]Y
*/

module horse_lights(
input [1:0]S,
input clk,
output reg [7:0]Y);

integer i;
reg sel;

always @(posedge clk)
	begin 
		Y[7:0]<=8'b00000000;
		sel<=0;
		if(S==2'b00)
		begin
			begin
				case(sel)
				0:
					begin
						for (i=0;i<2;i=i+1)
							begin 
								#1	Y[7:0]<=8'b10000000;
								#1	Y[7:0]<=8'b11000000;
								#1	Y[7:0]<=8'b11100000;
								#1	Y[7:0]<=8'b11110000;
								#1	Y[7:0]<=8'b11111000;
								#1	Y[7:0]<=8'b11111100;
								#1	Y[7:0]<=8'b11111110;
								#1	Y[7:0]<=8'b11111111;
								#1	Y[7:0]<=8'b01111111;
								#1	Y[7:0]<=8'b00111111;
								#1	Y[7:0]<=8'b00011111;
								#1	Y[7:0]<=8'b00001111;
								#1	Y[7:0]<=8'b00000111;
								#1	Y[7:0]<=8'b00000011;
								#1	Y[7:0]<=8'b00000001;
								#1	Y[7:0]<=8'b00000000;
							end 
								sel<=1;   
					end
				1:
					begin
						for (i=0;i<2;i=i+1)
							begin 
								#1	Y[7:0]<=8'b10000000;
								#1	Y[7:0]<=8'b11000000;
								#1	Y[7:0]<=8'b11100000;
								#1	Y[7:0]<=8'b11110000;
								#1	Y[7:0]<=8'b11111000;
								#1	Y[7:0]<=8'b11111100;
								#1	Y[7:0]<=8'b11111110;
								#1	Y[7:0]<=8'b11111111;
								#1	Y[7:0]<=8'b01111111;
								#1	Y[7:0]<=8'b00111111;
								#1	Y[7:0]<=8'b00011111;
								#1	Y[7:0]<=8'b00001111;
								#1	Y[7:0]<=8'b00000111;
								#1	Y[7:0]<=8'b00000011;
								#1	Y[7:0]<=8'b00000001;
								#1	Y[7:0]<=8'b00000000;

							end 
									S<=1;
					end	
			end	
		end		
	else if (S==2'b01)
		for (i=0;i<2;i=i+1)
		begin 
			#1	Y[7:0]<=8'b10000001;
			#1	Y[7:0]<=8'b11000011;
			#1	Y[7:0]<=8'b11100111;
			#1	Y[7:0]<=8'b11111111;
			#1	Y[7:0]<=8'b01111110;
			#1	Y[7:0]<=8'b00111100;
			#1	Y[7:0]<=8'b00011000;
			#1	Y[7:0]<=8'b00000000;
		end 
	else if (S==2'b10)
		for (i=0;i<2;i=i+1)
		begin 
			#1	Y[7:0]<=8'b11110001;
			#1	Y[7:0]<=8'b11110011;
			#1	Y[7:0]<=8'b11110111;
			#1	Y[7:0]<=8'b11111111;
			#1	Y[7:0]<=8'b11101111;
			#1	Y[7:0]<=8'b11001111;
			#1	Y[7:0]<=8'b10001111;
			#1	Y[7:0]<=8'b00001111;
			#1	Y[7:0]<=8'b11110000;
		end
	else 
		for (i=0;i<2;i=i+1)
		begin 
			#1	Y[7:0]<=8'b10000111;//分成两组灯，前四个灯为1组，后四个为2组，1组第1个灯亮，同时2组第1个灯不亮，第一组灯按从左到右依次点亮，之后按从左到右依次熄灭。然后第二组灯按同样的顺序依次熄灭与点亮；
			#1	Y[7:0]<=8'b11000011;
			#1	Y[7:0]<=8'b11100001;
			#1	Y[7:0]<=8'b11110000;
			#1	Y[7:0]<=8'b01111000;
			#1	Y[7:0]<=8'b00111100;
			#1	Y[7:0]<=8'b00011110;
			#1	Y[7:0]<=8'b00001111;
		end 
	end
		
endmodule




